library ieee;
use ieee.std_logic_1164.all;
entity G8BFA is
port(x,y : in std_logic_vector(7 downto 0);
Mgate : in std_logic;
cin : in std_logic;
sum : out std_logic_vector(7 downto 0);
cout : out std_logic);
end G8BFA;

architecture data1 of G8BFA is
signal cary : std_logic_vector(6 downto 0);


component GBFA is
port(A,B,Mgate,Cin : in std_logic;     
      Sout,Cout : out std_logic);    
end component;

begin 
a0 : GBFA port map (x(0),y(0),Mgate, cin,sum(0),cary(0));
a1 : GBFA port map (x(1),y(1),Mgate, cary(0),sum(1),cary(1));
a2 : GBFA port map (x(2), y(2),Mgate, cary(1), sum(2), cary(2));
a3 : GBFA port map (x(3), y(3),Mgate, cary(2), sum(3), cary(3));
a4 : GBFA port map (x(4), y(4),Mgate, cary(3), sum(4), cary(4));
a5 : GBFA port map (x(5), y(5),Mgate, cary(4), sum(5), cary(5));
a6 : GBFA port map (x(6), y(6),Mgate, cary(5), sum(6), cary(6));
a7 : GBFA port map (x(7), y(7),Mgate, cary(6), sum(7), cout);
end data1;
