library IEEE;
use IEEE.std_logic_1164.all;

entity GBFA is
port(A,B,Mgate,Cin : in std_logic;     
      Sout,Cout : out std_logic);    
end GBFA;

architecture struct of GBFA is
signal Ain: std_logic ;
component AND2 is
  port(P,Q : in std_logic;
        R : out std_logic);
end component;
component fa is
 port( X,Y,Z : in std_logic;
       U,V : out std_logic);
end component;
begin
a1:AND2 port map(A,Mgate,Ain);
a2:fa port map(Ain,B,Cin,Sout,Cout);
end struct;

