library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;

entity ALU is
port(A,B: in bit_vector(3 downto 0);
MS: in bit_vector(2 downto 0);
Ci: in bit;
S: out bit_vector(3 downto 0);
Co: out bit);
end ALU;

architecture structure of ALU is

component adder_4bit is
port(x,y : in bit_vector(3 downto 0);
cin : in bit;
sum : out bit_vector(3 downto 0);
cout : out bit);
end component;

signal t,u,v,w,o1,o2,p: bit_vector(3 downto 0);
signal t1,t2,t3,t4,n,o: bit;


begin
p<= NOT B;
n<='0';
o<= '1';
o1<= B"0000";
o2<= B"1111";
alu1: adder_4bit port map(A,B,Ci,sum=>t,cout=>t1); --Performing operation A + B + Cin
alu2: adder_4bit port map(A,p,o,sum=>u,cout=>t2);  --Performing operation A + B' + 1
alu3: adder_4bit port map(A,o1,o,sum=>v,cout=>t3); --Performing operation A + 1
alu4: adder_4bit port map(A,o2,n,sum=>w,cout=>t4);  -- Performing operationg A - 1 ( adding 2's compliment of 1 to A)
process(MS,t,u,v,w,t1,t2,t3,t4,n,o1)
begin
case MS is
when "000" =>
S<=t;
Co<=t1;
when "001" =>
S<=u;
Co<=t2;
when "010"=>
S<=v;
Co<=t3;
when "011"=>
S<=w;
Co<=t4;
when "100" =>  --Operation A
S <= A;
Co<=n;
when "101" =>  --Operation A and B
S <= A and B;
Co<=n;
when "110" =>  --Operation A or B
S <= A or B;
Co<=n;
when "111" =>  --Operation A'
S <= not A;
Co<=n;
when others =>
S <= o1;
Co<=n;
end case;
end process;
end structure;






